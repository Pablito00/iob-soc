assign gpio_input = 40;
